
//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 14-Jun-2024  1.0.0  DWW  Initial creation
// 13-Jul-2024  1.1.0  DWW  Added ability to fetch ABM data via DMA
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 1;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 13;
localparam VERSION_MONTH = 7;
localparam VERSION_YEAR  = 2024;

localparam RTL_TYPE      = 6142024;
localparam RTL_SUBTYPE   = 0;
